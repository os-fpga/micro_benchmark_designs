

module ram_inst_tdp_no_split_36 (
  input clock0, 
 //input clkA, clkB,
  input weA, weB,
  input [9:0] addrA, addrB,
  input [35:0] dinA, dinB, 
  output [35:0] doutA, doutB);


reg weA_reg, weB_reg;
reg [9:0]addrA_reg, addrB_reg;
reg [35:0] dinA_reg, dinB_reg;
reg [35:0]doutA, doutB;

wire [35 : 0]non_reg_doutA,non_reg_doutB;

always @(posedge clock0)
 begin
  weA_reg <= weA;
  weB_reg <= weB;
  addrA_reg <= addrA;
  addrB_reg <= addrB;
  dinA_reg <= dinA;
  dinB_reg <= dinB;
  doutA <= non_reg_doutA;
  doutB <= non_reg_doutB;
 end

parameter [80:0] MODE_BITS =81'hdb6;
// input clkA, clkB;
// input weA, weB;
// input [9:0] addrA, addrB;
// input [35:0] dinA, dinB;
// output [35:0] doutA, doutB;

 TDP36K  #(.MODE_BITS(81'hdb6))
  inst1(
    .ADDR_A1_i({ addrA_reg, 5'h00 }),
    .ADDR_A2_i({ addrA_reg[8:0], 5'h00 }),
    .ADDR_B1_i({ addrB_reg, 5'h00 }),
    .ADDR_B2_i({ addrB_reg[8:0], 5'h00 }),
    .BE_A1_i({1, 1}),
    .BE_A2_i({1, 1}),
    .BE_B1_i({1, 1}),
    .BE_B2_i({1, 1}),
    .CLK_A1_i(clock0),
    .CLK_A2_i(clock0),
    .CLK_B1_i(clock0),
    .CLK_B2_i(clock0),
    .FLUSH1_i(0),
    .FLUSH2_i(0),
    .RDATA_A1_o({non_reg_doutA[33:32],non_reg_doutA[15:0]}),
    .RDATA_A2_o({non_reg_doutA[35:34],non_reg_doutA[31:16]}),
    .RDATA_B1_o({non_reg_doutB[33:32],non_reg_doutB[15:0]}),
    .RDATA_B2_o({non_reg_doutB[35:34],non_reg_doutB[31:16]}),
    .REN_A1_i(),
    .REN_A2_i(),
    .REN_B1_i(),
    .REN_B2_i(),
    .RESET_ni(1),
    .WDATA_A1_i({dinA_reg[33:32],dinA_reg[15:0]}),
    .WDATA_A2_i({dinA_reg[35:34],dinA_reg[31:16]}),
    .WDATA_B1_i({dinB_reg[33:32],dinB_reg[15:0]}),
    .WDATA_B2_i({dinB_reg[35:34],dinB_reg[31:16]}),
    .WEN_A1_i(weA_reg),
    .WEN_A2_i(weA_reg),
    .WEN_B1_i(weB_reg),
    .WEN_B2_i(weB_reg)
  );
 

endmodule

/* Generated by Yosys 0.18+10 (git sha1 2b3815b19, gcc 9.4.0 -fPIC -Os) */

// (* top =  1  *)
// (* src = "/nfs_scratch/scratch/CompilerValidation/abdul_hameed/reggression/Compiler_Validation/RTL_testcases/Memory_Designs/Simple_dual_port_rams/ram_simple_dp_dc_512x32/rtl/ram_simple_dp_dc_512x32.v:1" *)
// module rams_sp_rwe(we, read_clock, write_clock, read_addr, write_addr, dout, din);
//   (* unused_bits = "32 33 34 35" *)
//   wire [35:0] \$auto$memory_bram.cc:844:replace_memory$48 ;
//   (* src = "/nfs_cadtools/raptor/instl_dir/bin/../share/yosys/rapidsilicon/genesis/brams_map.v:318.14-318.19" *)
//   (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35" *)
//   wire [35:0] \$techmap64\ram.0.0.0.DOBDO ;
//   (* src = "/nfs_scratch/scratch/CompilerValidation/abdul_hameed/reggression/Compiler_Validation/RTL_testcases/Memory_Designs/Simple_dual_port_rams/ram_simple_dp_dc_512x32/rtl/ram_simple_dp_dc_512x32.v:2" *)
//   input [31:0] din;
//   wire [31:0] din;
//   (* src = "/nfs_scratch/scratch/CompilerValidation/abdul_hameed/reggression/Compiler_Validation/RTL_testcases/Memory_Designs/Simple_dual_port_rams/ram_simple_dp_dc_512x32/rtl/ram_simple_dp_dc_512x32.v:5" *)
//   output [31:0] dout;
//   wire [31:0] dout;
//   (* src = "/nfs_scratch/scratch/CompilerValidation/abdul_hameed/reggression/Compiler_Validation/RTL_testcases/Memory_Designs/Simple_dual_port_rams/ram_simple_dp_dc_512x32/rtl/ram_simple_dp_dc_512x32.v:3" *)
//   input [8:0] read_addr;
//   wire [8:0] read_addr;
//   (* src = "/nfs_scratch/scratch/CompilerValidation/abdul_hameed/reggression/Compiler_Validation/RTL_testcases/Memory_Designs/Simple_dual_port_rams/ram_simple_dp_dc_512x32/rtl/ram_simple_dp_dc_512x32.v:4" *)
//   input read_clock;
//   wire read_clock;
//   (* src = "/nfs_scratch/scratch/CompilerValidation/abdul_hameed/reggression/Compiler_Validation/RTL_testcases/Memory_Designs/Simple_dual_port_rams/ram_simple_dp_dc_512x32/rtl/ram_simple_dp_dc_512x32.v:4" *)
//   input we;
//   wire we;
//   (* src = "/nfs_scratch/scratch/CompilerValidation/abdul_hameed/reggression/Compiler_Validation/RTL_testcases/Memory_Designs/Simple_dual_port_rams/ram_simple_dp_dc_512x32/rtl/ram_simple_dp_dc_512x32.v:3" *)
//   input [8:0] write_addr;
//   wire [8:0] write_addr;
//   (* src = "/nfs_scratch/scratch/CompilerValidation/abdul_hameed/reggression/Compiler_Validation/RTL_testcases/Memory_Designs/Simple_dual_port_rams/ram_simple_dp_dc_512x32/rtl/ram_simple_dp_dc_512x32.v:4" *)
//   input write_clock;
//   wire write_clock;
//   (* module_not_derived = 32'h00000001 *)
//   (* src = "/nfs_cadtools/raptor/instl_dir/bin/../share/yosys/rapidsilicon/genesis/brams_map.v:408.9-442.3" *)
//   TDP36K #(
//     .MODE_BITS(81'h00140281b6c0140140db6)
//   ) \ram.0.0.0  (
//     .ADDR_A1_i({ 1'h0, read_addr, 5'h00 }),
//     .ADDR_A2_i({ read_addr, 5'h00 }),
//     .ADDR_B1_i({ 1'h0, write_addr, 5'h00 }),
//     .ADDR_B2_i({ write_addr, 5'h00 }),
//     .BE_A1_i(2'h3),
//     .BE_A2_i(2'h3),
//     .BE_B1_i({ we, we }),
//     .BE_B2_i({ we, we }),
//     .CLK_A1_i(read_clock),
//     .CLK_A2_i(read_clock),
//     .CLK_B1_i(write_clock),
//     .CLK_B2_i(write_clock),
//     .FLUSH1_i(1'h0),
//     .FLUSH2_i(1'h0),
//     .RDATA_A1_o(dout[17:0]),
//     .RDATA_A2_o({ \$auto$memory_bram.cc:844:replace_memory$48 [35:32], dout[31:18] }),
//     .RDATA_B1_o(\$techmap64\ram.0.0.0.DOBDO [17:0]),
//     .RDATA_B2_o(\$techmap64\ram.0.0.0.DOBDO [35:18]),
//     .REN_A1_i(1'h1),
//     .REN_A2_i(1'h1),
//     .REN_B1_i(1'h0),
//     .REN_B2_i(1'h0),
//     .RESET_ni(1'h1),
//     .WDATA_A1_i(18'h3ffff),
//     .WDATA_A2_i(18'h3ffff),
//     .WDATA_B1_i(din[17:0]),
//     .WDATA_B2_i({ 4'hx, din[31:18] }),
//     .WEN_A1_i(1'h0),
//     .WEN_A2_i(1'h0),
//     .WEN_B1_i(we),
//     .WEN_B2_i(we)
//   );
//   assign \$auto$memory_bram.cc:844:replace_memory$48 [31:0] = dout;
// endmodule
